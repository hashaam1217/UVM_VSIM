`include "uvm_pkg.sv" 

